library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_ARITH.all;

entity imem is
    port(
        clk      : in  std_ulogic;
        addr     : in  std_ulogic_vector (6 downto 0);
        data     : out std_ulogic_vector (7 downto 0)
        );
end imem;
architecture BHV of imem is
    type ROM_TYPE is array (0 to 127) of std_ulogic_vector (7 downto 0);
    constant rom_content : ROM_TYPE := (
"10110000",    --IN R0
"00000000",    --NOP
"10110100",    --IN R1
"11011000",    --MOV R2, R0
"11011101",    --MOV R3, R1
"01000010",    --ADD R0, R2
"00000000",    --NOP
"00000000",    --NOP
"00000000",    --NOP
"00000000",    --NOP
"01000111",    --ADD R1, R3
"00000000",    --NOP
"00000000",    --NOP
"00000000",    --NOP
"11000000",    --OUT R0
"00000000",    --NOP
"00000000",    --NOP
"11000100",    --OUT R1
"00000000",    --NOP
"00000000",    --NOP
"11001000",    --OUT R2
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000");
begin
p1:    process (clk)
    variable add_in : integer := 0;
    begin
        if rising_edge(clk) then
            add_in := conv_integer(unsigned(addr));
            data <= rom_content(add_in);
        end if;
    end process;
end BHV;