library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_ARITH.all;


entity imem is
    port(
         clk      : in  std_ulogic;
         addr     : in  std_ulogic_vector (6 downto 0);
         data     : out std_ulogic_vector (7 downto 0)
         );
end imem;

architecture BHV of imem is

    type ROM_TYPE is array (0 to 127) of std_ulogic_vector (7 downto 0);

    constant rom_content : ROM_TYPE := (
  "00000000",	
  "10110000", -- input to r0 "11,0,0"
  "00000000",
	"11010100", -- move r0 to r1 "13,1,0"
  "00000000",
	"01000001", -- add r0, r1 "4,0,1"
  "00000000",
  "00000000",
  "00000000",
	"11000000", -- output r0 "12,0,0"
  "00000000",
  "00000000",
  "00000000",
  "00000000", 
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",	
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",	
	"00000000",	
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",	
	"00000000",	
	"00000000",
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",	
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",
	"00000000",
	"00000000",	
	"00000000",
	"00000000",
	"00000000",
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",
	"00000000",
	"00000000",	
	"00000000",
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",
	"00000000",
	"00000000",	
	"00000000",
	"00000000",
	"00000000",	
	"00000000",	
	"00000000",
	"00000000",
	"00000000",	
	"00000000",	
	"00000000",	
	"00000000",	
	"00000000",	
	"00000000",	
	"00000000",	
	"00000000",
	"00000000",	
	"00000000",	
	"00000000");
begin

p1:    process (clk)
	 variable add_in : integer := 0;
    begin
        if rising_edge(clk) then
					 add_in := conv_integer(unsigned(addr));
                data <= rom_content(add_in);
        end if;
    end process;
end BHV;
